* EESchema Netlist Version 1.1 (Spice format) creation date: 10/12/2012 17.55.44

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
D1  50 58 DIODE		
D2  61 58 DIODE		
CONN31  34 0 54 55 52 59 63 64 65 66 67 51 53 62 CONN_14		
CONN11  17 18 19 20 21 22 23 15 24 25 26 27 16 28 CONN_14		
CONN1  3 2 4 5 6 7 8 9 1 10 11 12 13 14 CONN_14		
CONN3  34 0 44 45 35 46 47 48 49 37 30 42 31 32 CONN_14		
XU1  36 29 BO2460		
XU3  38 39 SWITCH_DJ1235		
XU2  40 41 BO2460		
BAT1  34 42 JUMPER		
DIODE1  43 58 JUMPER		

.end
